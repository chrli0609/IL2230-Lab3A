module weight #(
    parameter N,
    parameter M,
    parameter WIDTH
)(
    //Need to have space for N*N*(M-1) memory segments
);

endmodule
