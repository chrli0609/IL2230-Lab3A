module data #() (


);

endmodule